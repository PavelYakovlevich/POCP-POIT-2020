----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:22:33 11/15/2020 
-- Design Name: 
-- Module Name:    lab4 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lab4 is
	 Generic (N : integer);
    Port ( DIN : in  STD_LOGIC_VECTOR (N-1 downto 0);
           DOUT : out  STD_LOGIC_VECTOR (N-1 downto 0);
           EN : in  STD_LOGIC);
end lab4;

architecture Behavioral of lab4 is

begin


end Behavioral;

