----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:57:57 10/25/2020 
-- Design Name: 
-- Module Name:    BI_STABLE_EL - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BI_STABLE_EL is
    Port ( I  : in   STD_LOGIC;
           Q  : out  STD_LOGIC;
           nQ : out  STD_LOGIC);
end BI_STABLE_EL;

architecture Behavioral of BI_STABLE_EL is

begin

	process (I)
	begin
		if I'event then
			Q  <= NOT(I);
			nQ <= I;
		end if;
	end process;

end Behavioral;

