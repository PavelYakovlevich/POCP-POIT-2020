----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:47:28 10/25/2020 
-- Design Name: 
-- Module Name:    DE_LATCH - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity DE_LATCH is
    Port ( D  : in   STD_LOGIC;
           E  : in   STD_LOGIC;
           Q  : out  STD_LOGIC;
           nQ : out  STD_LOGIC);
end DE_LATCH;

architecture Behavioral of DE_LATCH is

begin

	process(D, E)
	begin
		if E = '1' and (D = '1' or D = '0') then
			Q  <= D;
			nQ <= NOT(D);
		end if;
	end process;

end Behavioral;

