----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:23:28 09/29/2020 
-- Design Name: 
-- Module Name:    task4_1_demux - Structural 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity task4_1_demux is
    Port ( A : in  STD_LOGIC;
           S : in  STD_LOGIC;
           Z : out  STD_LOGIC;
           Z1 : out  STD_LOGIC);
end task4_1_demux;

architecture Structural of task4_1_demux is

begin



end Structural;

